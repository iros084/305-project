LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_ARITH.all;
USE  IEEE.STD_LOGIC_SIGNED.all;

entity start is
    port(pixel_row, pixel_col : in std_logic_vector(9 downto 0);
	       Clk, enable, mode_sel  : in std_logic;  -- if mode sel is '1', its game mode/ '0' is tutorial mode
         Red_out, Green_out, Blue_out : out std_logic);

end entity start;

architecture behaviour of start is

-- Signals for 2 digit counter
signal title_f_address : std_logic_vector(5 downto 0) := "000110";
signal title_l_address : std_logic_vector(5 downto 0) := "001100";
signal title_a_address : std_logic_vector(5 downto 0) := "000001";
signal title_p_address : std_logic_vector(5 downto 0) := "010000";
signal title_p1_address : std_logic_vector(5 downto 0) := "010000";
signal title_y_address : std_logic_vector(5 downto 0) := "011001";
signal title_b_address : std_logic_vector(5 downto 0) := "000010";
signal title_i_address : std_logic_vector(5 downto 0) := "001001";
signal title_r_address : std_logic_vector(5 downto 0) := "010010";
signal title_d_address : std_logic_vector(5 downto 0) := "000100";

signal play_p_address : std_logic_vector(5 downto 0) := "010000";
signal play_l_address : std_logic_vector(5 downto 0) := "001100";
signal play_a_address : std_logic_vector(5 downto 0) := "000001";
signal play_y_address : std_logic_vector(5 downto 0) := "011001";

signal tut_t_address : std_logic_vector(5 downto 0) := "010100";
signal tut_u_address : std_logic_vector(5 downto 0) := "010101";
signal tut_t1_address : std_logic_vector(5 downto 0) := "010100";
signal tut_o_address : std_logic_vector(5 downto 0) := "001111";
signal tut_r_address : std_logic_vector(5 downto 0) := "010010";
signal tut_i_address : std_logic_vector(5 downto 0) := "001001";
signal tut_a_address : std_logic_vector(5 downto 0) := "000001";
signal tut_l_address : std_logic_vector(5 downto 0) := "001100";

-- Signals for Sprite printing 
-- F L A P P Y B I R D
signal title_f_row : std_logic_vector(9 downto 0) := conv_std_logic_vector(120, 10);
signal title_f_col : std_logic_vector(9 downto 0) := conv_std_logic_vector(48, 10);
signal title_l_row : std_logic_vector(9 downto 0) := conv_std_logic_vector(120, 10);
signal title_l_col : std_logic_vector(9 downto 0) := conv_std_logic_vector(144, 10);
signal title_a_row : std_logic_vector(9 downto 0) := conv_std_logic_vector(120, 10);
signal title_a_col : std_logic_vector(9 downto 0) := conv_std_logic_vector(240, 10);
signal title_p_row : std_logic_vector(9 downto 0) := conv_std_logic_vector(120, 10);
signal title_p_col : std_logic_vector(9 downto 0) := conv_std_logic_vector(335, 10);
signal title_p1_row : std_logic_vector(9 downto 0) := conv_std_logic_vector(120, 10);
signal title_p1_col : std_logic_vector(9 downto 0) := conv_std_logic_vector(432, 10);
signal title_y_row : std_logic_vector(9 downto 0) := conv_std_logic_vector(120, 10);
signal title_y_col : std_logic_vector(9 downto 0) := conv_std_logic_vector(528, 10);
signal title_b_row : std_logic_vector(9 downto 0) := conv_std_logic_vector(200, 10);
signal title_b_col : std_logic_vector(9 downto 0) := conv_std_logic_vector(144, 10);
signal title_i_row : std_logic_vector(9 downto 0) := conv_std_logic_vector(200, 10);
signal title_i_col : std_logic_vector(9 downto 0) := conv_std_logic_vector(240, 10);
signal title_r_row : std_logic_vector(9 downto 0) := conv_std_logic_vector(200, 10);
signal title_r_col : std_logic_vector(9 downto 0) := conv_std_logic_vector(335, 10);
signal title_d_row : std_logic_vector(9 downto 0) := conv_std_logic_vector(200, 10);
signal title_d_col : std_logic_vector(9 downto 0) := conv_std_logic_vector(432, 10);


-- Flappy BIRD RGB
signal title_f_Red, title_f_Green, title_f_Blue,
       title_l_Red, title_l_Green, title_l_Blue,
       title_a_Red, title_a_Green, title_a_Blue,
       title_p_Red, title_p_Green, title_p_Blue,
       title_p1_Red, title_p1_Green, title_p1_Blue,
       title_y_Red, title_y_Green, title_y_Blue,
       title_b_Red, title_b_Green, title_b_Blue,
       title_i_Red, title_i_Green, title_i_Blue,
       title_r_Red, title_r_Green, title_r_Blue,
       title_d_Red, title_d_Green, title_d_Blue : std_logic;
            
signal Font_R : std_logic := '1';
Signal Font_G : std_logic := '1';
Signal Font_B : std_logic := '1';

Signal Font_Multiplier : integer := 4;
signal select_multiplier : integer := 3;

component Sprite_Printer is	
  port(pixel_row, pixel_col, anchor_row, anchor_col : in std_logic_vector(9 downto 0);
       sprite_red, sprite_green, sprite_blue : in std_logic;
       multiplier : in integer range 1 to 4;
       address : in std_logic_vector (5 downto 0);
       enable, clk : in std_logic;
       red_out, green_out, blue_out : out std_logic);
end component Sprite_printer;

	begin
          title_f: sprite_printer port map(pixel_row, pixel_col, title_f_row, title_f_col, Font_R, Font_G, Font_B, Font_Multiplier, title_f_address, enable, CLK, title_f_Red, title_f_Green, title_f_Blue);
	  title_l: sprite_printer port map(pixel_row, pixel_col, title_l_row, title_l_col, Font_R, Font_G, Font_B, Font_Multiplier, title_l_address, enable, CLK, title_l_Red, title_l_Green, title_l_Blue);
	  title_a: sprite_printer port map(pixel_row, pixel_col, title_a_row, title_a_col, Font_R, Font_G, Font_B, Font_Multiplier, title_a_address, enable, CLK, title_a_Red, title_a_Green, title_a_Blue);
	  title_p: sprite_printer port map(pixel_row, pixel_col, title_p_row, title_p_col, Font_R, Font_G, Font_B, Font_Multiplier, title_p_address, enable, CLK, title_p_Red, title_p_Green, title_p_Blue);
 	  title_p1: sprite_printer port map(pixel_row, pixel_col, title_p1_row, title_p1_col, Font_R, Font_G, Font_B, Font_Multiplier, title_p1_address, enable, CLK, title_p1_Red, title_p1_Green, title_p1_Blue);
	  title_y: sprite_printer port map(pixel_row, pixel_col, title_y_row, title_y_col, Font_R, Font_G, Font_B, Font_Multiplier, title_y_address, enable, CLK, title_y_Red, title_y_Green, title_y_Blue);
	  title_b: sprite_printer port map(pixel_row, pixel_col, title_b_row, title_b_col, Font_R, Font_G, Font_B, Font_Multiplier, title_b_address, enable, CLK, title_b_Red, title_b_Green, title_b_Blue);
	  title_i: sprite_printer port map(pixel_row, pixel_col, title_i_row, title_i_col, Font_R, Font_G, Font_B, Font_Multiplier, title_i_address, enable, CLK, title_i_Red, title_i_Green, title_i_Blue);
	  title_r: sprite_printer port map(pixel_row, pixel_col, title_r_row, title_r_col, Font_R, Font_G, Font_B, Font_Multiplier, title_r_address, enable, CLK, title_r_Red, title_r_Green, title_r_Blue);
	  title_d: sprite_printer port map(pixel_row, pixel_col, title_d_row, title_d_col, Font_R, Font_G, Font_B, Font_Multiplier, title_d_address, enable, CLK, title_d_Red, title_d_Green, title_d_Blue);
	
	
    play_RED <= not(mode_sel);
    tut_RED <= mode_sel;
	  
    Red_out <= title_f_R_out and title_l_R_out and title_a_R_out and title_p_R_out and title_p1_R_out and title_y_R_out and title_b_R_out and title_i_R_out and title_r_R_out and title_d_R_out; 
    Green_out <= title_f_G_out and title_l_G_out and title_a_G_out and title_p_G_out and title_p1_G_out and title_y_G_out and title_b_G_out and title_i_G_out and title_r_G_out and title_d_G_out; 
    Blue_out <= title_f_B_out and title_l_B_out and title_a_B_out and title_p_B_out and title_p1_B_out and title_y_B_out and title_b_B_out and title_i_B_out and title_r_B_out and title_d_B_out; 
end architecture;